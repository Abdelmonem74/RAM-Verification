package classes_pack;
    `include "transaction.svh"
    `include "sequencer.svh"
    `include "driver.svh"
    `include "monitor.svh"
    `include "subscriber.svh"
    `include "scoreboard.svh"
    `include "env.svh"
endpackage