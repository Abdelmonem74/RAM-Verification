package pack1;
    import uvm_pkg::*;
    import config_pack::*;
    `include "uvm_macros.svh";
    `include "my_sequence_item.svh"
    `include "my_sequence.svh"
    `include "my_sequencer.svh"
    `include "my_driver.svh"
    `include "my_monitor.svh"
    `include "my_scoreboard.svh"
    `include "my_subscriber.svh"
    `include "my_agent.svh"
    `include "my_env.svh"
    `include "my_test.svh"

    
endpackage
