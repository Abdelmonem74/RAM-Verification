module top ();

    import uvm_pkg::*;
    import pack1::*;
    import config_pack::*;

    ////////////////////////////////////////////////////////////////////////////////////////////////////////
    //////////////////////////////////////////    CLOCK      ///////////////////////////////////////////
    ////////////////////////////////////////////////////////////////////////////////////////////////////////
    bit clk_tb;

    ////////////////////////////////////////////////////////////////////////////////////////////////////////
    ///////////////////////////////////////   INTERFACE INSTANT  ///////////////////////////////////////////
    ////////////////////////////////////////////////////////////////////////////////////////////////////////
    intf ram_cif();

    ////////////////////////////////////////////////////////////////////////////////////////////////////////
    ///////////////////////////////////////     DUT INSTANCE     ///////////////////////////////////////////
    ////////////////////////////////////////////////////////////////////////////////////////////////////////
    ram  dut (.intf1(ram_cif.dut)); 
    //virtual intf.tb vif;

    ////////////////////////////////////////////////////////////////////////////////////////////////////////
    ///////////////////////////////////////    CLOCK GENERATOR   ///////////////////////////////////////////
    ////////////////////////////////////////////////////////////////////////////////////////////////////////
    assign ram_cif.clk = clk_tb;
    always #(clk_period/2) clk_tb = ~clk_tb;

    initial begin
        uvm_config_db #(virtual intf)::set(null, "uvm_test_top", "my_vif",ram_cif);
        $display("run_test!!!!!!");
        run_test("my_test");
        
    end
endmodule