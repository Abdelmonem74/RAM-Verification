package config_pack;
    parameter int ADDR_WIDTH = 4;
    parameter int DATA_WIDTH = 32;
    parameter int clk_period = 10;

endpackage