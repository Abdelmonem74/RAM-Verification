`timescale 1ps/1ps
module tbench ();
////////////////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////    CLOCK      ///////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////////
bit clk_tb;
////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////   PACKAGE IMPORTION   ///////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////////
import classes_pack::*;
import config_pack::*;

////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////   INTERFACE INSTANT  ///////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////////
intf  ram_cif();
virtual intf.tb class_vif;

////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////   ENVIRONMENT CLASS  ///////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////////
env env1;
////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////     DUT INSTANCE     ///////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////////
ram  dut (.intf1(ram_cif.dut)); 

////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////    CLOCK GENERATOR   ///////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////////
assign ram_cif.clk = clk_tb;
always #(clk_period/2) clk_tb = ~clk_tb;


initial begin
////////////////////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////    Connecting vif with cif   //////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////////
    class_vif = ram_cif.tb;

////////////////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////    ENVIRONMENT CLASS   //////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////////
    env1 = new(class_vif);
////////////////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////   TestCases   //////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////////
    env1.run();
    
    env1.end_sim();
end
endmodule